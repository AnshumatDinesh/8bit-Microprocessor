module Control_Unit (
    input[]
);
    
endmodule