module Decoder_8bit (
    input wire [7:0] I,
    output reg [255:0]O
);
    
endmodule